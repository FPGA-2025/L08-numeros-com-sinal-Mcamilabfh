module numeros_com_sinal(
    input signed [7:0] entrada_signed_1,
    input signed [3:0] entrada_signed_2,
    input [7:0] entrada_unsigned_1,
    input [3:0] entrada_unsigned_2,
    input [1:0] codigo,
    output reg [7:0] saida
);

always @(*) begin
    case (codigo)
        2'b00: saida = entrada_signed_1 + entrada_signed_2;  // signed + signed
        2'b01: saida = entrada_unsigned_1 + entrada_unsigned_2; // unsigned + unsigned
        2'b10: saida = entrada_unsigned_1 + entrada_signed_1; // unsigned + signed
        2'b11: saida = entrada_unsigned_1 + entrada_signed_2; // unsigned + signed
        default: saida = 8'b0; // Só pra garantir uma saída padrão
    endcase
    end

endmodule